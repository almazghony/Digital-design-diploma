module bcd(input i0, i1, i2, i3, i4, i5, i6, i7, i8, i9,
            output reg o0, o1, o2, o3);
    always @(*) begin
        case ({i0, i1, i2, i3, i4, i4, i5, i6, i7, i8, i9})
            'b0000000001 : {o0, o1, o2, o3} = 'b0000;
            'b0000000010 : {o0, o1, o2, o3} = 'b0001;
            'b0000000100 : {o0, o1, o2, o3} = 'b0010;
            'b0000001000 : {o0, o1, o2, o3} = 'b0011;
            'b0000010000 : {o0, o1, o2, o3} = 'b0100;
            'b0000100000 : {o0, o1, o2, o3} = 'b0101;
            'b0001000000 : {o0, o1, o2, o3} = 'b0110;
            'b0010000000 : {o0, o1, o2, o3} = 'b0111;
            'b0100000000 : {o0, o1, o2, o3} = 'b1000;
            'b1000000000 : {o0, o1, o2, o3} = 'b1001;
            

        endcase
    end 
endmodule